module ALU(
    input wire clk,
    input wire rst_n,
    input wire [7:0] A,
    input wire [7:0] B,
    input wire start,
    input wire [2:0] opcode,
    output wire [15:0] result,
    output wire done
);


endmodule: ALU