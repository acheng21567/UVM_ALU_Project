typedef uvm_sequencer#(sequence_item) sequencer;